module TOP();
   flashloader i1 (.noe_in(1'd0));
endmodule
